// Chris Kenyon and Brandon Nguyen
// CPU Test bench

`timescale 1ns / 100ps

module CPU_tb;
  reg clk, reset;
  wire[31:0] instruction, dataOut, dataIn, instructionAddress, dataAddress;
  wire MemRead, MemWrite;
  
Memory memory(instructionAddress, instruction, dataAddress, dataIn, MemRead, MemWrite, dataOut);  
CPU cpu(reset, instructionAddress, instruction, dataAddress, dataIn, MemRead, MemWrite, dataOut, clk);

initial begin
  reset = 0;
  clk = 0;
  reset = 1;
  #5
  reset = 0;
end

always
  #10 clk = !clk;

always #100 $display("R0: %h R1: %h \n", cpu.regFile.regFile[0], cpu.regFile.regFile[1]);
  always #100 $display("R2: %h R3: %h \n", cpu.regFile.regFile[2], cpu.regFile.regFile[3]);
  always #100 $display("R4: %h R5: %h \n", cpu.regFile.regFile[4], cpu.regFile.regFile[5]);
  always #100 $display("R6: %h R7: %h \n", cpu.regFile.regFile[6], cpu.regFile.regFile[7]);
  always #100 $display("R8: %h R9: %h \n", cpu.regFile.regFile[8], cpu.regFile.regFile[9]);
  always #100 $display("R100: %h R11: %h \n", cpu.regFile.regFile[100], cpu.regFile.regFile[11]);
  always #100 $display("R12: %h R13: %h \n", cpu.regFile.regFile[12], cpu.regFile.regFile[13]);
  always #100 $display("R14: %h R15: %h \n", cpu.regFile.regFile[14], cpu.regFile.regFile[15]);
  always #100 $display("R16: %h R17: %h \n", cpu.regFile.regFile[16], cpu.regFile.regFile[17]);
  always #100 $display("R18: %h R19: %h \n", cpu.regFile.regFile[18], cpu.regFile.regFile[19]);
  always #100 $display("R20: %h R21: %h \n", cpu.regFile.regFile[20], cpu.regFile.regFile[21]);
  always #100 $display("R22: %h R23: %h \n", cpu.regFile.regFile[22], cpu.regFile.regFile[23]);
  always #100 $display("R24: %h R25: %h \n", cpu.regFile.regFile[24], cpu.regFile.regFile[25]);
  always #100 $display("R26: %h R27: %h \n", cpu.regFile.regFile[26], cpu.regFile.regFile[27]);
  always #100 $display("R28: %h R29: %h \n", cpu.regFile.regFile[28], cpu.regFile.regFile[29]);
  always #100 $display("R30: %h R31: %h \n", cpu.regFile.regFile[30], cpu.regFile.regFile[31]);

endmodule
